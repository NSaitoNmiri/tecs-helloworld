import (<sPrint.cdl>);

celltype tOutput {
	entry sPrint ePrint;
};

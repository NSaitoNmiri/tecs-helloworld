signature sPrint {
	void print([in, string] const char *str);
};
